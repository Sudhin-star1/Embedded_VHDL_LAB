LIBRARY ieee;

USE ieee.std_logic_1164.ALL;

ENTITY HA_tb IS

END HA_tb;

ARCHITECTURE behavior OF HA_tb IS 

    COMPONENT Half_Adder

    PORT(

         A : IN  std_logic;

         B : IN  std_logic;

         S : OUT  std_logic;

         C : OUT  std_logic

        );

    END COMPONENT;


   signal A : std_logic := '0';

   signal B : std_logic := '0';


   signal S : std_logic;

   signal C : std_logic;


BEGIN


   uut: Half_Adder PORT MAP (

          A => A,

          B => B,

          S => S,

          C => C

        );



   stim_proc: process

   begin		


      wait for 100 ns;	

		

	 A <= '0';

    B <= '0';

    wait for 10 ns;

	 

    A <= '0';

    B <= '1';

    wait for 10 ns;

	 

    A <= '1';

    B <= '0';

    wait for 10 ns;

	 

    A <= '1';

    B <= '1';

    wait for 10 ns;


      wait;

   end process;



END;